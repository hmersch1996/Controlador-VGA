library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Driver_VGA is
    Port ( CLK : in  STD_LOGIC;
           REINICIO : in  STD_LOGIC;
           HSYNC : out  STD_LOGIC;
           VSYNC : out  STD_LOGIC;
			  SELECTOR: in STD_LOGIC;
			  
           Red : out  STD_LOGIC_VECTOR (2 downto 0);
			  Green : out  STD_LOGIC_VECTOR (2 downto 0);
			  Blue : out  STD_LOGIC_VECTOR (2 downto 0)
);
end Driver_VGA;

  architecture Behavioral of Driver_VGA is

signal CLK50: STD_LOGIC :='0';
signal CLK25: STD_LOGIC :='0';

constant HD: integer := 639; -- 639 DISPLAY HORIZONTAL (640)
constant HFP: integer := 16; --  16 BORDE DERECHO (porche frontal)
constant HSP: integer := 96; --  96 SYNC PULSE (sincronizacion horizontal)
constant HBP: integer := 48; --  48 BORDE IZQUIERDO (porche trasero)

constant VD: integer := 479; -- 479 DISPLAY VERTICAL(480) 
constant VFP: integer := 10; --  10 RIGHT BORDER (porche frontal)
constant VSP: integer := 2;  --   2 SYNC PULSE (sincronizacion vertical)
constant VBP: integer := 33; --  33 LEFT BORDER (porche trasero)

type mem is array (160 downto 0) of std_logic_vector(159 downto 0);
type mem2 is array (63 downto 0) of std_logic_vector(319 downto 0);

signal Matriz : mem;
signal MatrizL : mem2;

signal hpos: integer :=0;
signal vpos: integer :=0;

signal videoOn: STD_LOGIC :='0';
begin

MatrizL(0) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(1) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(2) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(3) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(4) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(5) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(6) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(7) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(8) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(9) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(10) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(11) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(12) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(13) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(14) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(15) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111110000000000111111111111111111111111111";
MatrizL(16) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111100000000111111111111111111111111111111";
MatrizL(17) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111100000001111111111111111111111111111111";
MatrizL(18) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111100000011111111111111111111111111111111";
MatrizL(19) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111000000011111111111111111111111111111111";
MatrizL(20) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111000000011111111111111111111111111111111";
MatrizL(21) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111110000000011111111111111111111111111111111";
MatrizL(22) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010011111111111111111110000010011111111111111111111111111111111";
MatrizL(23) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010001111111111111111100000110011111111111111111111111111111111";
MatrizL(24) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111110000011001111111111111111100000110011111111111111111111111111111111";
MatrizL(25) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111110000011000111111111111111000000110011111111111111111111111111111111";
MatrizL(26) <= "11111111111111111111111111111111111100000001111111111111111000000111111111111111001111111111111111000001111100011111111111111100000001111111111100001111000111111111111100000111111111111000000011111111111111100000011111111111111111100000011111111111111110000011100111111111111111000001110011111111111111111111111111111111";
MatrizL(27) <= "11111111111111111111111111111111110000000000011111111111100000000001111111111111000001111111111100000000011100000111111111110000000000011111111000000011000001111100000000000011111111100000000000111111111110000000000111111111111110000000000111111111111110000011100011111111111110000001110011111111111111111111111111111111";
MatrizL(28) <= "11111111111111111111111111111111100000111100001111111111000001111000011111111111000000011111111100000000001100000000111111100000111100000111111000000001000000011100000000000001111111000001111000011111111000000111100001111111111100000111110001111111111110000011110011111111111110000011110011111111111111111111111111111111";
MatrizL(29) <= "11111111111111111111111111111111000001111110000111111110000011111110001111111111000000001111111000001111100100000000111111000001111111000011111100011100000000001111111000001111111110000011111100001111111000001111111000111111111000001111111000111111111110000011110011111111111110000011110011111111111111111111111111111111";
MatrizL(30) <= "11111111111111111111111111111111000011111111000011111100000111111110000111111111000001111111111000011111110000000111111110000011111111100011111111111110000001111111111000001111111110000111111110000111110000011111111000011111110000011111111100011111111110000011111001111111111100000111110011111111111111111111111111111111";
MatrizL(31) <= "11111111111111111111111111111111000011111111000011111100000111111111000111111111000001111111111000011111111100000111111100000111111111110001111111111111000001111111111100001111111110000111111110000111110000011111111100011111110000011111111110011111111110000011111001111111111100000111110011111111111111111111111111111111";
MatrizL(32) <= "11111111111111111111111111111111000011111111000011111100000111111111000011111111000011111111110000011111111100000111111100000111111111110000111111111111000001111111111100001111111110000111111110000111110000011111111100001111100000111111111110001111111110000011111000111111111000001111110011111111111111111111111111111111";
MatrizL(33) <= "11111111111111111111111111111111000011111111000011111110001111111111100011111111000011111111110000011111111100000111111000001111111111110000111111111111000001111111111100001111111110000111111110000111111000111111111110001111100000111111111110001111111110000011111100111111111000001111110011111111111111111111111111111111";
MatrizL(34) <= "11111111111111111111111111111111000011111111100111111111111111111111100001111111000011111111110000011111111100000111111000001111111111110000111111111111000001111111111100001111111110000111111111001111111111111111111110000111100000000000000000000111111110000011111100011111110000011111110011111111111111111111111111111111";
MatrizL(35) <= "11111111111111111111111111111111000001111111111111111111111111111111100001111111000011111111110000011111111100000111111000001111111111110000011111111111000001111111111100001111111110000011111111111111111111111111111110000111100000000000000000000111111110000011111110011111110000011111110011111111111111111111111111111111";
MatrizL(36) <= "11111111111111111111111111111111000000001111111111111111111111111111100001111111000011111111110000011111111100000111110000011111111111110000011111111111000001111111111100001111111110000000011111111111111111111111111110000111111111111111111110000111111110000011111110001111100000011111110011111111111111111111111111111111";
MatrizL(37) <= "11111111111111111111111111111111000010000011111111111111111111111111100001111111000011111111110000011111111100000111110000011111111111110000011111111111000001111111111100001111111110000100000111111111111111111111111110000111111111111111111110000111111110000011111111001111100000111111110011111111111111111111111111111111";
MatrizL(38) <= "11111111111111111111111111111111000011110000111111111111111111111111100001111111000011111111110000011111111100000111110000011111111111110000011111111111000001111111111100001111111110000111100001111111111111111111111110000111111111111111111110000111111110000011111111000111000000111111110011111111111111111111111111111111";
MatrizL(39) <= "11111111111111111111111111111111000011111100001111111111111111111111100001111111000011111111110000011111111100000111111000011111111111110000011111111111000001111111111100001111111110000111111000011111111111111111111110000111111111111111111110000111111110000011111111100111000001111111110011111111111111111111111111111111";
MatrizL(40) <= "11111111111111111111111111111111000011111110000111111111111111111111000001111111000011111111110000011111111100000111111000011111111111110000011111111111000001111111111100001111111110000111111100001111111111111111111100000111111111111111111110000111111110000011111111100010000001111111110011111111111111111111111111111111";
MatrizL(41) <= "11111111111111111111111111111111000011111111000011111011111111111111000001111111000001111111110000011111111100000111111000011111111111110000011111111111000001111111111000001111111110000111111110000111101111111111111100000111101111111111111100000111111110000011111111110010000011111111110011111111111111111111111111111111";
MatrizL(42) <= "11111111111111111111111111111111000011111111100001111001111111111111000001111111000001111111110000011111111100000111111000011111111111110000011111111111000001111111111100001111111110000111111110000111110111111111111100000111101111111111111100000111111110000011111111110000000011111111110011111111111111111111111111111111";
MatrizL(43) <= "11111111111111111111111111111111000011111111100001111101111111111110000011111111000011111111110000011111111100000111111000011111111111100000111111111111000001111111111000001111111110000111111111000011110111111111111000001111100111111111111000001111111110000011111111111000000111111111110011111111111111111111111111111111";
MatrizL(44) <= "11111111111111111111111111111111000011111111100001111100111111111100000011111111000011111111110000011111111100000111111100001111111111100000111111111111000001111111111000001111111110000111111111000011110011111111110000001111110011111111110000001111111110000011111111111000000111111111110011111111111111111111111111111111";
MatrizL(45) <= "11111111111111111111111111111111000011111111000001111110011111111000000011111111000011111111110000011111111100000111111110001111111111000001111111111111000001111111111000001111111110000111111111000011111001111111100000001111110011111111100000011111111110000011111111111000001111111111110011111111111111111111111111111111";
MatrizL(46) <= "11111111111111111111111111111110000001111111000001111110000111110000000111111111000001111111110000011111111100000111111110001111111111000001111111111111000001111011111000001111111110000011111110000011111000011111000000011111111000111111000000011111111110000011111111111100001111111111110011111111111111111111111111111111";
MatrizL(47) <= "11111111111111111111111111110110000000011110000001111111000000000000001111111111000001111111110000011111111100000111111111000111111110000011111111111111000001111100110000001111101100000000111100000011111100000000000000111111111100000000000000111111111110000011111111111100011111111111100001111111111111111111111111111111";
MatrizL(48) <= "11111111111111111111111111111000000011000000000011111111100000000000011111111110000000111111100000001111111000000011111111100001111000000111111111111110000000111110000000011111110000000110000000000111111110000000000001111111111110000000000001111111111000000000111111111110011111111111000000111111111111111111111111111111";
MatrizL(49) <= "11111111111111111111111111111100000111100000000111111111110000000000111111110000000000001110000000000001100000000000111111110000000000001111111111110000000000001110000000111111111000000111000000001111111111000000000011111111111111000000000011111111000000000000000111111110111111111000000000000111111111111111111111111111";
MatrizL(50) <= "11111111111111111111111111111110000111111000001111111111111110000011111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111100001111111111100001111110000011111111111110000001111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(51) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(52) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(53) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(54) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(55) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(56) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(57) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(58) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(59) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(60) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(61) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(62) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
MatrizL(63) <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";

Matriz(0) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(1) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(2) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(3) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(4) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(5) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(6) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(7) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(8) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(9) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(10) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(11) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(12) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(13) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(14) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(15) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(16) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(17) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(18) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(19) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(20) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(21) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(22) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(23) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(24) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(25) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(26) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(27) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(28) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(29) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(30) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(31) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(32) <= "0000000000000000000000000000000000000000000000000000000000000000000000000010011010010011000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(33) <= "0000000000000000000000000000000000000000000000000000000000000000000000010110010010010001100010000000000000000000000000000000000000000000000000000000000000000000";
Matriz(34) <= "0000000000000000000000000000000000000000000000000000000000000000001100010110010001010000100111000000000000000000000000000000000000000000000000000000000000000000";
Matriz(35) <= "0000000000000000000000000000000000000000000000000000000000000011001010011000010010010000101101001000000000000000000000000000000000000000000000000000000000000000";
Matriz(36) <= "0000000000000000000000000000000000000000000000000000000000000001001111011001011110010001001111001001000000000000000000000000000000000000000000000000000000000000";
Matriz(37) <= "0000000000000000000000000000000000000000000000000000000000000001001001000000000000000010010001010111000000000000000000000000000000000000000000000000000000000000";
Matriz(38) <= "0000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000001011001000000000000000000000000000000000000000000000000000000000000";
Matriz(39) <= "0000000000000000000000000000000000000000000000000000001100000001100000000001111111111000000000010010000000000000000000000000000000000000000000000000000000000000";
Matriz(40) <= "0000000000000000000000000000000000000000000000000000010010000010000000100000000000000000010000000010000001110000000000000000000000000000000000000000000000000000";
Matriz(41) <= "0000000000000000000000000000000000000000000000000000010011000000000000000000000000000000000011000000000010011000000000000000000000000000000000000000000000000000";
Matriz(42) <= "0000000000000000000000000000000000000000000000000110010001000000100000000000000000000000000000010000000100010000000000000000000000000000000000000000000000000000";
Matriz(43) <= "0000000000000000000000000000000000000000000000001001001110000010000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000";
Matriz(44) <= "0000000000000000000000000000000000000000000000000011100000001000000000000000000000000000000000000001000011100011000000000000000000000000000000000000000000000000";
Matriz(45) <= "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010001001101000000000000000000000000000000000000000000000000";
Matriz(46) <= "0000000000000000000000000000000000000000000000000000100000000000000000000011111111111000000000000000001000011101000000000000000000000000000000000000000000000000";
Matriz(47) <= "0000000000000000000000000000000000000000000000000001000100000000000000111111111111111111110000000000000010000010000000000000000000000000000000000000000000000000";
Matriz(48) <= "0000000000000000000000000000000000000000000000000000000000000000000111111111001100100111111100000000000001000010011100000000000000000000000000000000000000000000";
Matriz(49) <= "0000000000000000000000000000000000000000001110000000000000000000011110011111001100100110010111100000000000100000100010000000000000000000000000000000000000000000";
Matriz(50) <= "0000000000000000000000000000000000000000001101110000000000000001111010011001001100000110000011111000000000010000100110000000000000000000000000000000000000000000";
Matriz(51) <= "0000000000000000000000000000000000000000000111000000000000000011110010011001001100000000000011011100000000001000101100000000000000000000000000000000000000000000";
Matriz(52) <= "0000000000000000000000000000000000000000000010000000000000001110111111111001000000000000010000001111000000000100011001100000000000000000000000000000000000000000";
Matriz(53) <= "0000000000000000000000000000000000000001110011000000000000011100111001011001000000100000010000001001100000000010000110000000000000000000000000000000000000000000";
Matriz(54) <= "0000000000000000000000000000000000000001010000000000000000111100100001011001000000100001000001000001110000000001001100001000000000000000000000000000000000000000";
Matriz(55) <= "0000000000000000000000000000000000000000010010000000000001100101001011111001000000000100010000100000111000000000000011101000000000000000000000000000000000000000";
Matriz(56) <= "0000000000000000000000000000000000000000011100000000000011100101011111111001100000000000001100010000001100000000000010111000000000000000000000000000000000000000";
Matriz(57) <= "0000000000000000000000000000000000000011000000000000000101100110110000011011000000000000000010001000000110000000010010000000000000000000000000000000000000000000";
Matriz(58) <= "0000000000000000000000000000000000000000100000000000001101110111101001111011000110000111100001100100000011000000000001000110000000000000000000000000000000000000";
Matriz(59) <= "0000000000000000000000000000000000000000010000000000011101011111100011111011000111000100011100010110100001100000001000001000000000000000000000000000000000000000";
Matriz(60) <= "0000000000000000000000000000000000001100010000000000111110011111111100011111000111000000000111001010100000110000000100001001000000000000000000000000000000000000";
Matriz(61) <= "0000000000000000000000000000000000000011100000000000111110011111100000011111000011000000000011100101000000110000000000000110000000000000000000000000000000000000";
Matriz(62) <= "0000000000000000000000000000000000010000000000000001101100010010111111111111000000000100000000111011010000111000000000011000000000000000000000000000000000000000";
Matriz(63) <= "0000000000000000000000000000000000011110000000000011001101100010110110011011000000000100000000011101010010011000000000000000100000000000000000000000000000000000";
Matriz(64) <= "0000000000000000000000000000000000001000000000000011001101000011111111011010000000000000000000001110100011001100000000001010000000000000000000000000000000000000";
Matriz(65) <= "0000000000000000000000000000000000000100000000000111001101010100011110011110000000000000000000000011001011000100000001001001110000000000000000000000000000000000";
Matriz(66) <= "0000000000000000000000000000000000011100000000000111001101101100111010011110000000000000000000010001101010000110000000001111000000000000000000000000000000000000";
Matriz(67) <= "0000000000000000000000000000000000000000000000001101101111110001110010011111111111100000000000001000111010000110000000100000010000000000000000000000000000000000";
Matriz(68) <= "0000000000000000000000000000000000111000000000001111111111111110110010011100000000000000010000000100010010010010000000100000100000000000000000000000000000000000";
Matriz(69) <= "0000000000000000000000000000000001001100000000001011111111111100110010011100000000000000010000000010000110000011000000000011000000000000000000000000000000000000";
Matriz(70) <= "0000000000000000000000000000000010000100000000011010011001101100110010011111110000010000010000000001000110000011000000000011111000000000000000000000000000000000";
Matriz(71) <= "0000000000000000000000000000000000000100000000011010001001111110110010010000010000000000010010000000100100101011100000010000000000000000000000000000000000000000";
Matriz(72) <= "0000000000000000000000000000000000000000000000011010000001000100110010110000110000010000000010000000010010101011100000010000000000000000000000000000000000000000";
Matriz(73) <= "0000000000000000000000000000000011111000000000011010110001001100110010100000110000011000000010000011011010001010100000000011111000000000000000000000000000000000";
Matriz(74) <= "0000000000000000000000000000000000000000000000011010010101001100110011100000110000011100000010000111101000001010100000000000000000000000000000000000000000000000";
Matriz(75) <= "0000000000000000000000000000000001100000000000111011010101011100110011000000110000001100000010000000100100011010100000000000001000000000000000000000000000000000";
Matriz(76) <= "0000000000000000000000000000000011011000000000111001101110110100110011000000110000001110000010000000110100011010100000000001100000000000000000000000000000000000";
Matriz(77) <= "0000000000000000000000000000000000001000000000111011111111100100110110000000110000001111000010000000010110010010110000000000110000000000000000000000000000000000";
Matriz(78) <= "0000000000000000000000000000000000001000000000111011011111100100110110000001110000000111000000000001010010010000110000000000001000000000000000000000000000000000";
Matriz(79) <= "0000000000000000000000000000000011110000000000111011001101111100111100000000110000000111100000000011111000110000110000000001111100000000000000000000000000000000";
Matriz(80) <= "0000000000000000000000000000000000000000000000111111011011111100111100000000110000000111110000000011101000110000110000000000000000000000000000000000000000000000";
Matriz(81) <= "0000000000000000000000000000000000000000000000111101110011101100111000001000110000000011110000000000101000100000110000000000111000000000000000000000000000000000";
Matriz(82) <= "0000000000000000000000000000000011100000000000111100010001001100111000001000110000000010111000000000100101100100110000000001000000000000000000000000000000000000";
Matriz(83) <= "0000000000000000000000000000000001000000000000111100010001001100110000001100000000000000010100000000100101100100110000000010000000000000000000000000000000000000";
Matriz(84) <= "0000000000000000000000000000000000010000000000011100010001001100110000001100000000000000100000000000110101001000100000000001000000000000000000000000000000000000";
Matriz(85) <= "0000000000000000000000000000000011111000000000011010110101001101100100000100000000000001000000000000110001011000100000000000111100000000000000000000000000000000";
Matriz(86) <= "0000000000000000000000000000000000000000000000011011010101011101100000000011111111110000000000000000110000110000100000000000000000000000000000000000000000000000";
Matriz(87) <= "0000000000000000000000000000000000000000000000011011101001111111000000000000000000000000000000000000100001100011100000010000000000000000000000000000000000000000";
Matriz(88) <= "0000000000000000000000000000000000000000000000011011111111101111110000000000000000000000000000000000100011100011100000010000000000000000000000000000000000000000";
Matriz(89) <= "0000000000000000000000000000000000000000000000011001011111101111111001000000000000000000000000000000100111000010000000000000000000000000000000000000000000000000";
Matriz(90) <= "0000000000000000000000000000000000000000000000001001001111111010111111100000000000000000011000000000100110011011000000000000000000000000000000000000000000000000";
Matriz(91) <= "0000000000000000000000000000000000000000000000001001001100110010110011110000000000000000011000000010101100111011000000000000000000000000000000000000000000000000";
Matriz(92) <= "0000000000000000000000000000000000000000000000001111111100010001110010110001100000011000010000000010011001000010000000100000000000000000000000000000000000000000";
Matriz(93) <= "0000000000000000000000000000000000001000000000000111111110001001110011111001111000111100010000000100110100000110000000000001000000000000000000000000000000000000";
Matriz(94) <= "0000000000000000000000000000000000001100000000000111100010000101111010011001111100111100010000000101101000100110000000000011000000000000000000000000000000000000";
Matriz(95) <= "0000000000000000000000000000000000000000000000000011100000010101111110011000011100100110000010001010010000110100000000000000000000000000000000000000000000000000";
Matriz(96) <= "0000000000000000000000000000000000000000000000000011110011000111111110011001001100100110000100000100100000011000000000000000000000000000000000000000000000000000";
Matriz(97) <= "0000000000000000000000000000000000000000000000000001111000101110110011011001001100100110000100001000000000011000000000000000000000000000000000000000000000000000";
Matriz(98) <= "0000000000000000000000000000000000000000000000000001101110011111110001111001001100100110000000010000000000110000000000000000000000000000000000000000000000000000";
Matriz(99) <= "0000000000000000000000000000000000000000000000000000111111111110011000111001001100100110000001000000010000110000000000000000000100000000000000000000000000000000";
Matriz(100) <= "0000000000000000000000000000000000000000000000000000011101100110000110111111001100101111000010000001100001100000000000100000000000000000000000000000000000000000";
Matriz(101) <= "0000000000000000000000000000000000000001111000000000001101100111000001011111111111111111100000000110000011000000000001011000001000000000000000000000000000000000";
Matriz(102) <= "0000000000000000000000000000000000000111001000000000001101111110100100111111111111111111100000000000000110000000000001011100000000000000000000000000000000000000";
Matriz(103) <= "0000000000000000000000000000000000000000110000000000000111110000010001111111111111111111100000000000000100000000000000010000010000000000000000000000000000000000";
Matriz(104) <= "0000000000000000000000000000000000000000100000000000000011101000111111111111111111111111100000000000011100000000000000000000000000000000000000000000000000000000";
Matriz(105) <= "0000000000000000000000000000000000000001000100000000000001111110000001111111111111111111100000000001110000000000000101100000100000000000000000000000000000000000";
Matriz(106) <= "0000000000000000000000000000000000000000011000000000000000011111111110011111111101111111110000000011100000000000000110100000000000000000000000000000000000000000";
Matriz(107) <= "0000000000000000000000000000000000000000010001100000000000001110110010011111111101111111010011001111000000000000000011000001000000000000000000000000000000000000";
Matriz(108) <= "0000000000000000000000000000000000000000000010010000000000000111110010011111111100111111010011011100000000000000010001000000000000000000000000000000000000000000";
Matriz(109) <= "0000000000000000000000000000000000000000001111110000000000000001111010011011111100111110010011111000000000000001101101000000000000000000000000000000000000000000";
Matriz(110) <= "0000000000000000000000000000000000000000000001000100000000000000011110011001001100100110010111100000000000000000000100000100000000000000000000000000000000000000";
Matriz(111) <= "0000000000000000000000000000000000000000000010000010000000000000000111111001001100100110111110000000000000000010000100001000000000000000000000000000000000000000";
Matriz(112) <= "0000000000000000000000000000000000000000000000001110000000000000000000111111111111111111110000000000000000000001000100000000000000000000000000000000000000000000";
Matriz(113) <= "0000000000000000000000000000000000000000000001001100100000000000000000000011111111111100000000000000000000010001100000000000000000000000000000000000000000000000";
Matriz(114) <= "0000000000000000000000000000000000000000000000111001000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000";
Matriz(115) <= "0000000000000000000000000000000000000000000000010010010000000000000000000101011000101100000000000000000000100100100000000000000000000000000000000000000000000000";
Matriz(116) <= "0000000000000000000000000000000000000000000000000100100010000000000000000101011001100100000000000000000000110011000000000000000000000000000000000000000000000000";
Matriz(117) <= "0000000000000000000000000000000000000000000010000000111110000000000000000100011001100100000000000000011000010000000000000000000000000000000000000000000000000000";
Matriz(118) <= "0000000000000000000000000000000000000000000000000001100100010000000000000000000000000100000000000000101000001000000000000000000000000000000000000000000000000000";
Matriz(119) <= "0000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000010000100010000000000000000000000000000000000000000000000000000";
Matriz(120) <= "0000000000000000000000000000000000000000000000000000001000110001000000000000000000000000000000000111000100000000000000000000000000000000000000000000000000000000";
Matriz(121) <= "0000000000000000000000000000000000000000000000000000000010010000100000000000000000000000000001100101100010000000000000000000000000000000000000000000000000000000";
Matriz(122) <= "0000000000000000000000000000000000000000000000000010000001100100100000100000000000000000000110100111110000000000000000000000000000000000000000000000000000000000";
Matriz(123) <= "0000000000000000000000000000000000000000000000000000000000001000101011101000001110011100000100010110000000000000000000000000000000000000000000000000000000000000";
Matriz(124) <= "0000000000000000000000000000000000000000000000000000010000000111001110001000000010110000000110010010000000000000000000000000000000000000000000000000000000000000";
Matriz(125) <= "0000000000000000000000000000000000000000000000000000000100000000001001001000000110100010000011110000000000000000000000000000000000000000000000000000000000000000";
Matriz(126) <= "0000000000000000000000000000000000000000000000000000000000000000000001001000000010100010000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(127) <= "0000000000000000000000000000000000000000000000000000000000010000000000000000000010011110000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(128) <= "0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(129) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(130) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(131) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(132) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(133) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(134) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(135) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(136) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(137) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(138) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(139) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(140) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(141) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(142) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(143) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(144) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(145) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(146) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(147) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(148) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(149) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(150) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(151) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(152) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(153) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(154) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(155) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(156) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(157) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(158) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
Matriz(159) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

--Como es necesario trabajar con un reloj de 25 MHz, es necesario crearlo a partir del reloj de 100 MHz.
--Esta funcion nos permite obtener un reloj de 50 MHz. 
--Solo cuando el reloj de 100 MHz llega a un flanco positivo, el reloj de 50 MHz cambia de estado
divisor_de_clock:process(CLK)
begin
	if(CLK'event and CLK='1') then 
		CLK50 <= NOT CLK50;
	end if;
end process;

--Esta funcion nos permite obtener un reloj de 50 MHz. 
--Solo cuando el reloj de 50 MHz llega a un flanco positivo, el reloj de 25 MHz cambia de estado
divisor_de_clock50:process(CLK50)
begin
	if(CLK50'event and CLK50='1') then
		CLK25 <= NOT CLK25;
	end if;
end process;

--Aqui se realiza el conteo de la posicion horizontal.
contador_posicion_horizontal:process(CLK25,REINICIO)
begin
	if(REINICIO='1') then --Si el reinicio se activa, hpos se resetea
		hpos <=0;
	elsif(CLK25'event and CLK25='1') then
		if (hpos=(HD+HFP+HSP+HBP)) then --Si hpos llega a la ultima posicion posible, se reinicia
			hpos <=0;
		else
			hpos <= hpos+1;
		end if;
	end if;
end process;

--Aqui se realiza el conteo de la posicion vertical.
contador_posicion_vertical:process(CLK25,REINICIO,hpos)
begin
	if(REINICIO='1') then 							--Si el reinicio se activa, vpos se resetea
		vpos <=0;
	elsif(CLK25'event and CLK25='1') then
		if (hpos=(HD+HFP+HSP+HBP)) then 			--vpos cambia cuando hpos llega a su posicion final
			if (vpos=(VD+VFP+VSP+VBP)) then 		--si vpos llega a su posicion final, vpos se resetea
				vpos <=0;
			else
				vpos <= vpos+1;
			end if;
		end if;
	end if;
end process;

--Aqui se realiza la sincronizacion horizontal
sincronizacion_horizontal:process(CLK25,REINICIO,hpos)
begin
	if(REINICIO='1') then											--Si el reinicio se activa, HSYNC se resetea
		HSYNC <= '0';
	elsif(CLK25'event and CLK25='1') then
		if ((hpos <= (HD+HFP)) or (hpos>HD+HFP+HSP)) then  --Si hpos esta entre el porche delantero y trasero, HSYNC se activa
			HSYNC <='1';
		else
			HSYNC <='0';
		end if;
	end if;
end process;

--Aqui se realiza la sincronizacion vertical
sincronizacion_vertical:process(CLK25,REINICIO,vpos)
begin
	if(REINICIO='1') then                                 --Si el reinicio se activa, VSYNC se resetea
		VSYNC <= '0';
	elsif(CLK25'event and CLK25='1') then
		if ((vpos <= (VD+VFP)) or (Vpos>VD+VFP+VSP)) then  --Si vpos esta entre el porche delantero y trasero, VSYNC se activa
			VSYNC <='1';
		else
			VSYNC <='0';
		end if;
	end if;
end process;

--Aqui definimos si se muestra o no algo en pantalla
video_on:process(CLK25,REINICIO, hpos,vpos)
begin
	if(REINICIO='1') then										--Si el reinicio se activa, videoON se resetea
		videoON <= '0';
	elsif(CLK25'event and CLK25='1') then
		if (hpos <=HD and vpos <=VD) then					--Si hpos y vpos estan dentro del rango visible, el video se activa
			videoON <= '1';
		else
			videoON <= '0';
		end if;
	end if;
end process;


draw: process (VideoON,REINICIO, hpos, vpos)   
variable offset : natural;
variable offset2 : natural;
variable xint, yint : integer;
variable color : std_logic;
begin  
--Escalado horizontal y horizontal
xint := hpos/2; 
yint := vpos/4; 
	if(REINICIO = '1')then --Se verifica si el reset esta activo
		Red <= "000"; -- Se asigna loa tonos a los colores Rojo, Verde y Azul
		Green <= "000"; 
		Blue <= "000"; 
	elsif(CLK25'event and CLK25='1') then 
		if videoON = '1' then 
			--Se modifica el offset que queda de la imagen luego del escalado
			offset := ( yint * 120)+( xint ); 
			offset2 := (xint * 240 ) + (yint);
			--Se controla la imagen a mostrar
			if selector='1' then 
				--Se determina el rango de la imagen 1
				if (hpos>=0 and hpos<640) AND (vpos>160 and vpos<320) then 
						--Se guarda cada bit de la imagen para luego asignarle el respectivo color
						color := MatrizL(yint-220)(xint); 
						Red <= "000";
						Green <= "000"; 
						Blue <= (others=>color);
				end if;
				
			else --Se selecciona la otra imagen a mostrar
				color := Matriz(yint-240)(xint-100);
					Red <="111";
					Green <=(others=>color);
					Blue <=(others=>color);
			end if;
			--En caso que no haya imagen a visualizar en cierto sector, se le asigna este color
			else 
			Red <="000";
			Green <="000";
			Blue <="000";
		end if;
	end if;
end process;

 
end Behavioral;



